--Kushal Kumar Gupta 2020CS10355

library IEEE;
use IEEE.std_logic_1164.all;

entity do_nothing is
	--does nothing
end do_nothing;

architecture no_arch of do_nothing is
begin
	--does nothing
end no_arch;